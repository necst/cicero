`timescale 1ns/1ps

package basic_block_task_package;

   

endpackage : basic_block_task_package 