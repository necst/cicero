
package basic_block_task_package;

   

endpackage : basic_block_task_package 