`timescale 1ns / 10ps

import instruction::*;

module regex_cpu_pipelined_split_tb();
    parameter CLOCK_SEMI_PERIOD = 5  ;

    parameter  PC_WIDTH          = 8;
    parameter  CHARACTER_WIDTH   = 8;
    parameter  MEMORY_WIDTH      = 16;
    parameter  MEMORY_ADDR_WIDTH = 11;

    logic                             clk                               ;
    logic                             reset                             ; 
    logic[CHARACTER_WIDTH-1:0]        current_character                 ;
    logic                             input_pc_valid                    ;
    logic[PC_WIDTH-1:0]               input_pc                          ;
    logic                             input_pc_ready                    ;
    logic                             memory_ready                      ;
    logic[MEMORY_ADDR_WIDTH-1:0]      memory_addr                       ;
    logic[MEMORY_WIDTH-1     :0]      memory_data                       ;
    logic                             memory_valid                      ;
    logic                             output_pc_is_directed_to_current  ;
    logic                             output_pc_valid                   ;
    logic[PC_WIDTH-1:0]               output_pc                         ;
    logic                             output_pc_ready                   ;
    logic                             accepts                           ;
    logic                             running                           ;

    regex_cpu_pipelined #(
        .PC_WIDTH             (PC_WIDTH             ),
        .CHARACTER_WIDTH      (CHARACTER_WIDTH      ),
        .MEMORY_WIDTH         (MEMORY_WIDTH         ),
        .MEMORY_ADDR_WIDTH    (MEMORY_ADDR_WIDTH    ),
        .FIFO_WIDTH_POWER_OF_2(2                    )   
    )a_cpu_under_test(
        .clk                               ( clk                               ),
        .reset                             ( reset                             ), 
        .current_character                 ( current_character                 ),
        .input_pc_valid                    ( input_pc_valid                    ),
        .input_pc                          ( input_pc                          ), 
        .input_pc_ready                    ( input_pc_ready                    ),
        .memory_ready                      ( memory_ready                      ),
        .memory_addr                       ( memory_addr                       ),
        .memory_data                       ( memory_data                       ),
        .memory_valid                      ( memory_valid                      ),
        .output_pc_is_directed_to_current  ( output_pc_is_directed_to_current  ),
        .output_pc_valid                   ( output_pc_valid                   ),
        .output_pc                         ( output_pc                         ),
        .output_pc_ready                   ( output_pc_ready                   ),
        .accepts                           ( accepts                           ),
        .running                           ( running                           )
);

    // clock generator  
    always begin
        #CLOCK_SEMI_PERIOD clk = ~ clk;
    end

    task load_pc_and_supply_memory(  input reg[PC_WIDTH-1    :0] pc,
                                    input reg[MEMORY_WIDTH-1     :0] value
                                    );
    begin
        
        input_pc_valid <= 1'b1;
        input_pc       <= pc;
        @(posedge clk);
        memory_ready   <= 1'b1;
        @(posedge clk);
        input_pc_valid <= 1'b0;
        memory_data  <= value;
        memory_ready <= 1'b0;
        if(memory_valid !== 1'b1)
        begin
            $display("regex_cpu does not wait memory");
            $stop();
        end
        if(memory_addr !== pc)
        begin
            $display("regex_cpu address mismatch %h != %h", memory_addr, pc);
            $stop();
        end
        @(posedge clk);
        if(running !== 1'b1)
        begin
            $display("regex_cpu seems not having received instruction");
            $stop();
        end
        if(memory_valid == 1'b1)
        begin
            $display("regex_cpu want something frem memory even if it had just fetched!");
            $stop();
        end
        
    end
    endtask

    task wait_2pc_unordered_output(
                        input reg[MEMORY_ADDR_WIDTH-1:0]expected0_pc,
                        input reg                       expected0_is_directed_to_current,
                        input reg[MEMORY_ADDR_WIDTH-1:0]expected1_pc,
                        input reg                       expected1_is_directed_to_current
                        );
    begin
        logic zero_ok=1'b0;
        logic one_ok=1'b0;
        while(output_pc_valid == 1'b0 )
            @(posedge clk);
            if(~running)
            begin
                $display("regex_cpu stopped running without producing any pc!");
                $stop();
            end
        repeat(2)
            begin
            @(posedge clk);
            output_pc_ready    <= 1'b1;

            if( output_pc_valid !== 1'b1)
            begin
                $display("regex_cpu didn't need to produce pc!");
                $stop();
            end
            if(output_pc == expected0_pc)
            begin 
                if(output_pc_is_directed_to_current !== expected0_is_directed_to_current)
                begin
                    $display("regex_cpu is directed to current %h != %h", output_pc_is_directed_to_current, expected0_is_directed_to_current);
                    $stop();
                end
                else
                begin
                    zero_ok=1'b1;
                end
            end
            else if(output_pc == expected1_pc)
            begin 
                if(output_pc_is_directed_to_current !== expected1_is_directed_to_current)
                begin
                    $display("regex_cpu is directed to current %h != %h", output_pc_is_directed_to_current, expected1_is_directed_to_current);
                    $stop();
                end
                else
                begin
                    zero_ok=1'b1;
                end
            end
            else
            begin
                $display("regex_cpu output pc %h not in [ %h, %h] ", output_pc, expected0_pc, expected1_pc);
                $stop();
            end
            @(posedge clk);
            output_pc_ready    <=1'b0;
        end
        @(posedge clk);
        if(running)
        begin
            $display("regex_cpu still has work to do!");
            $stop();
        end
        
        
    end
    endtask



    initial begin
        reg [PC_WIDTH-1:0] a_pc, another_pc;
        reg [PC_WIDTH-1:0] max_pc, max_another_pc;
        
        max_pc          = 64;
        max_another_pc  = 64; 
        
        input_pc_valid  = 1'b0;
        memory_ready    = 1'b0;
        output_pc_ready = 1'b0;
        clk             = 1'b0;
        reset          <= 1'b0;
        @(posedge clk);
        reset          <= 1'b1;
        @(posedge clk);
        reset          <= 1'b0;
        repeat(30) @(posedge clk);

        for ( a_pc = 0 ; a_pc < max_pc ; a_pc+=1 ) begin
            for(another_pc = 0 ; another_pc < max_another_pc; another_pc+=1)begin
                current_character <= 8'h00;
                
                load_pc_and_supply_memory(a_pc,{SPLIT,another_pc });
                wait_2pc_unordered_output(a_pc+8'h01, 1'b1, another_pc, 1'b1);
                $display("OK %h -> %h,%h", a_pc, a_pc+1, another_pc);
                
                repeat (10)
                    begin
                        @(posedge clk);
                        if( output_pc_valid == 1'b1)
                        begin
                            $display("regex_cpu didn't need to produce pc!");
                            $stop();
                        end
                        if( running == 1'b1)
                        begin
                            $display("regex_cpu still working");
                            $stop();
                        end
                    end
            end
        end
        

        $display("OK");
        $finish();

    end

endmodule